LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
USE IEEE.math_real.all;

ENTITY Memory IS
    GENERIC ( n : INTEGER := 16; m : INTEGER := 20);     
    PORT (
        EXT_CLK         	: IN  STD_LOGIC;
        EXT_INTR		: IN  STD_LOGIC;

	IR1_IN				: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	IR2_IN				: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	PC	      		: IN  STD_LOGIC_VECTOR(31 DOWNTO 0); 
	SP	      	    	: IN  STD_LOGIC_VECTOR(31 DOWNTO 0);

------------------------------------------------------------------------------
	
	Rsrc1			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	Rdst1			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);

	Read_Enable1		: IN  STD_LOGIC;
	Write_Enable1		: IN  STD_LOGIC;
	ALU_As_Address1		: IN  STD_LOGIC;
	SP_As_Address1		: IN  STD_LOGIC;
	PC_As_Data1 		: IN  STD_LOGIC;

	ALU1_OUT		: IN  STD_LOGIC_VECTOR( 31 DOWNTO 0);

-------------------------------------------------------------------------------	

	Rsrc2			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	Rdst2			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);

	Read_Enable2		: IN  STD_LOGIC;
	Write_Enable2		: IN  STD_LOGIC;
	ALU_As_Address2		: IN  STD_LOGIC;
	SP_As_Address2		: IN  STD_LOGIC;
	PC_As_Data2 		: IN  STD_LOGIC;
	
	ALU2_OUT		: IN  STD_LOGIC_VECTOR( 31 DOWNTO 0);

	RET1_OUT			: OUT STD_LOGIC;
	RET2_OUT			: OUT STD_LOGIC;
	Memory_OUT		: OUT STD_LOGIC_VECTOR( 31 DOWNTO 0)  
    );
END ENTITY;

ARCHITECTURE arch_Memory OF Memory IS

SIGNAL mem_address   : STD_LOGIC_VECTOR(m-1 DOWNTO 0);
SIGNAL mem_read	     : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL mem_data	     : STD_LOGIC_VECTOR(31 DOWNTO 0);

SIGNAL mem_PC_data   : STD_LOGIC;
SIGNAL Read_Enable   : STD_LOGIC;
SIGNAL Write_Enable  : STD_LOGIC;
SIGNAL SP_Address    : STD_LOGIC;

SIGNAL ZERO_VECTOR   : STD_LOGIC_VECTOR(15 DOWNTO 0) := (others => '0');

BEGIN
						  -- both wont be 1 at the same time (Hazard)
Read_Enable  <= Read_Enable1 or Read_Enable2;     -- if Ch1 or Ch2 wants to read
Write_Enable <= Write_Enable1 or Write_Enable2;   -- If Ch1 or Ch2 wants to write
mem_PC_data  <= PC_As_Data1 or PC_As_Data2;
SP_Address   <= SP_As_Address1 or SP_As_Address2;

Data_Memory:
ENTITY work.memory_data
GENERIC MAP(n => 16, m => 20)
PORT MAP(
	CLK       => EXT_CLK,
	RD        => Read_Enable,
	WR        => Write_Enable,
	PC_Data   => mem_PC_data,
	Address   => mem_address,
	WriteData => mem_data,
	
	ReadData  => mem_read
);



	
	mem_address <= SP(m-1 DOWNTO 0) when SP_Address = '1' and (Read_Enable = '1' or Write_Enable = '1') -- PUSH Instruction
		else ALU1_OUT(m-1 DOWNTO 0) when ALU_As_Address1 = '1' and (Read_Enable = '1' or Write_Enable = '1') -- pop instruction Ch1 --> take ALU 1 out
		else ALU2_OUT(m-1 DOWNTO 0) when ALU_As_Address2 = '1' and (Read_Enable = '1' or Write_Enable = '1') -- pop instruction Ch2 --> take ALU 2 out
		else ZERO_VECTOR(3 DOWNTO 0) & Rsrc1 when ALU_As_Address1 = '0' and Read_Enable1 = '1'  -- Load Instruction
		else ZERO_VECTOR(3 DOWNTO 0) & Rsrc2 when ALU_As_Address2 = '0' and Read_Enable2 ='1' 
		else ZERO_VECTOR(3 DOWNTO 0) & Rdst1 when SP_Address = '0' and Write_Enable1 = '1'  -- store instruction
		else ZERO_VECTOR(3 DOWNTO 0) & Rdst2 when SP_Address = '0' and Write_Enable2 = '1'; 


	mem_data <= std_logic_vector(unsigned(PC)+1) when mem_PC_data = '1' and Write_Enable = '1' -- Call instruction -- *****NOTE PC or PC+1  not sure yet
		else ZERO_VECTOR(15 downto 0) & Rdst1 when SP_As_Address1 = '1' and Write_Enable = '1' -- Push instruction in Ch1  *** May change it to Rsrc not Rdst
		else ZERO_VECTOR(15 downto 0) & Rdst2 when SP_As_Address2 = '1' and Write_Enable = '1'	-- Push Instruction in Ch2  *** Same as above
		else ZERO_VECTOR(15 downto 0) & Rsrc1 when Write_Enable1 = '1' and Write_Enable = '1' -- Store instruction in Ch1
		else ZERO_VECTOR(15 downto 0) & Rsrc2 when Write_Enable2 = '1' and Write_Enable = '1';

	RET1_OUT <= '1' when IR1_IN(15 DOWNTO 10) = "100110"
				else '0';
	RET2_OUT <= '1' when IR2_IN(15 DOWNTO 10) = "100110"
				else '0';
	
	Memory_OUT <= mem_read;


END ARCHITECTURE;