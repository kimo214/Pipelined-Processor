LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
USE IEEE.math_real.all;

ENTITY Memory IS
    GENERIC ( n : INTEGER := 16; m : INTEGER := 10);     
    PORT (
        EXT_CLK         	: IN  STD_LOGIC;
        EXT_INTR		: IN  STD_LOGIC;
	EXT_RST			: IN  STD_LOGIC; 

	PC	      		: IN  STD_LOGIC_VECTOR(31 DOWNTO 0); 
	SP	      	    	: IN  STD_LOGIC_VECTOR(31 DOWNTO 0);

------------------------------------------------------------------------------
	
	Rsrc1			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	Rdst1			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);

	Read_Enable1		: IN  STD_LOGIC;
	Write_Enable1		: IN  STD_LOGIC;
	ALU_As_Address1		: IN  STD_LOGIC;
	SP_As_Address1		: IN  STD_LOGIC;
	PC_As_Data1 		: IN  STD_LOGIC;

	ALU1_OUT		: IN  STD_LOGIC_VECTOR( 31 DOWNTO 0);

-------------------------------------------------------------------------------	

	Rsrc2			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	Rdst2			: IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);

	Read_Enable2		: IN  STD_LOGIC;
	Write_Enable2		: IN  STD_LOGIC;
	ALU_As_Address2		: IN  STD_LOGIC;
	SP_As_Address2		: IN  STD_LOGIC;
	PC_As_Data2 		: IN  STD_LOGIC;
	
	ALU2_OUT		: IN  STD_LOGIC_VECTOR( 31 DOWNTO 0);


	Memory_OUT		: OUT STD_LOGIC_VECTOR( 31 DOWNTO 0)  
    );
END ENTITY;

ARCHITECTURE arch_Memory OF Memory IS

SIGNAL mem_address   : STD_LOGIC_VECTOR(m-1 DOWNTO 0);
SIGNAL mem_read	     : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL mem_data	     : STD_LOGIC_VECTOR(31 DOWNTO 0);

SIGNAL mem_PC_data   : STD_LOGIC;
SIGNAL Read_Enable   : STD_LOGIC;
SIGNAL Write_Enable  : STD_LOGIC;
SIGNAL SP_Address    : STD_LOGIC;

SIGNAL ZERO_VECTOR   : STD_LOGIC_VECTOR(15 DOWNTO 0) := (others => '0');

BEGIN
						  -- both wont be 1 at the same time (Hazard)
Read_Enable  <= Read_Enable1 or Read_Enable2;     -- if Ch1 or Ch2 wants to read
Write_Enable <= Write_Enable1 or Write_Enable2;   -- If Ch1 or Ch2 wants to write
mem_PC_data  <= PC_As_Data1 or PC_As_Data2;
SP_Address   <= SP_As_Address1 or SP_As_Address2;

Data_Memory:
ENTITY work.memory_data
GENERIC MAP(n => 16, m => 10)
PORT MAP(
	CLK       => EXT_CLK,
	RD        => Read_Enable,
	WR        => Write_Enable,
	PC_Data   => mem_PC_data,
	Address   => mem_address,
	WriteData => mem_data,
	
	ReadData  => mem_read
);


PROCESS(EXT_CLK, Read_Enable, Write_Enable)
BEGIN
	IF(Read_Enable = '1' or Write_Enable = '1') THEN
		-- Determine Which address to use
		IF(SP_Address = '1') THEN  					-- PUSH Instruction
			mem_address <= SP;
		ELSIF(ALU_As_Address1 = '1') THEN			-- pop instruction Ch1 --> take ALU 1 out
			mem_address <= ALU1_OUT;
		ELSIF(ALU_As_Address2 = '1') THEN			-- pop instruction Ch2 --> take ALU 2 out
			mem_address <= ALU2_OUT;
		ELSIF(Read_Enable1 = '1') THEN				-- Load Instruction
			mem_address <= ZERO_VECTOR & Rsrc1;
		ELSIF(Read_Enable2 ='1') THEN
			mem_address <= ZERO_VECTOR & Rsrc2;
		ELSIF(Write_Enable1 = '1') THEN				-- store instruction
			mem_address <= ZERO_VECTOR & Rdst1;
		ELSIF(Write_Enable2 = '1') THEN
			mem_address <= ZERO_VECTOR & Rdst2;
		END IF;

		IF(Write_Enable = '1') THEN
			IF(mem_PC_data = '1') THEN           	 -- Call instruction
				mem_data <= PC;               	 	 -- *****NOTE PC or PC+1  not sure yet
			ELSIF(SP_As_Address1 = '1') THEN     	 -- Push instruction in Ch1  *** May change it to Rsrc not Rdst
				mem_data <= Rdst1;	
			ELSIF(SP_As_Address2 = '1') THEN     	 -- Push Instruction in Ch2  *** Same as above
				mem_data <= Rdst2; 
			ELSIF(Write_Enable1 = '1') THEN      	 -- Store instruction in Ch1
				mem_data <= Rsrc1;
			ELSIF(Write_Enable2 = '1') THEN      	 -- Store instruction in Ch2
				mem_data <= Rsrc2;
			END IF;
		END IF;

		IF(Read_Enable = '1' and Rising_Edge(EXT_CLK)) THEN
			Memory_OUT <= mem_read;
		END IF;
	END IF;
END PROCESS;

END ARCHITECTURE;